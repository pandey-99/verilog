
 `timescale 1ns/1ps
 module test;
  reg [3:0] A,B;
  reg Cin;
  wire [3:0] S;
  wire Cout;
 
    full_adder uut(.A(A),.B(B),.Cin(Cin),.S(S),.Cout(Cout));
   initial  begin

    A=4'b0000;
    B=4'b0000;
    Cin=1'b0;
    
  
    
    $dumpfile("full_adder_tb.vcd");
    $dumpvars(0,test);
     
    #10 A=4'b0000; B=4'b0001;Cin=0;
    #10 A=4'b0000; B=4'b0010;
    #10 A=4'b0000; B=4'b0011;
    #10 A=4'b0000; B=4'b0100;
    #10 A=4'b0000; B=4'b0101;
    #10 A=4'b0000; B=4'b0110;
    #10 A=4'b0000; B=4'b0111;
    #10 A=4'b0000; B=4'b1000;
    #10 A=4'b0000; B=4'b1001;
    #10 A=4'b0000; B=4'b1010;
    #10 A=4'b0000; B=4'b1011;
    #10 A=4'b0000; B=4'b1100;
    #10 A=4'b0000; B=4'b1101;   
    #10 A=4'b0000; B=4'b1111;
    #10 A=4'b0001; B=4'b0010;
    #10 A=4'b0010; B=4'b0011;
    #10 A=4'b0011; B=4'b0100;
    #10 A=4'b0100; B=4'b0101;
    #10 A=4'b0101; B=4'b0110;
    #10 A=4'b0110; B=4'b0111;
    #10 A=4'b0111; B=4'b1000;
    #10 A=4'b1000; B=4'b1001;
    #10 A=4'b1001; B=4'b1010;
    #10 A=4'b1010; B=4'b1010;
    #10 A=4'b1011; B=4'b1011;
    #10 A=4'b1110; B=4'b1100;
    #10 A=4'b1111; B=4'b1101;   
    #10 A=4'b1101; B=4'b1111;
    #10 A=4'b0000; B=4'b0000;Cin=1;
    #10 A=4'b0000; B=4'b0010;
    #10 A=4'b0000; B=4'b0011;
    #10 A=4'b0000; B=4'b0100;
    #10 A=4'b0000; B=4'b0101;
    #10 A=4'b0000; B=4'b0110;
    #10 A=4'b0000; B=4'b0111;
    #10 A=4'b0000; B=4'b1000;
    #10 A=4'b0000; B=4'b1001;
    #10 A=4'b0000; B=4'b1010;
    #10 A=4'b0000; B=4'b1011;
    #10 A=4'b0000; B=4'b1100;
    #10 A=4'b0000; B=4'b1101;   
    #10 A=4'b0000; B=4'b1111;
    #10 A=4'b0001; B=4'b0010;
    #10 A=4'b0010; B=4'b0011;
    #10 A=4'b0011; B=4'b0100;
    #10 A=4'b0100; B=4'b0101;
    #10 A=4'b0101; B=4'b0110;
    #10 A=4'b0110; B=4'b0111;
    #10 A=4'b0111; B=4'b1000;
    #10 A=4'b1000; B=4'b1001;
    #10 A=4'b1001; B=4'b1010;
    #10 A=4'b1010; B=4'b1010;
    #10 A=4'b1011; B=4'b1011;
    #10 A=4'b1110; B=4'b1100;
    #10 A=4'b1111; B=4'b1101;   
    #10 A=4'b1101; B=4'b1111;
    #10 $finish;
  end
endmodule
